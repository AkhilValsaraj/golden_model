`define BR	0000
`define ADD	0001
`define LD	0010
`define ST	0011
`define JSR	0100	//JSRR
`define AND	0101
`define LDR	0110
`define STR	0111
`define RTI	1000
`define NOT	1001
`define LDI	1010
`define STI	1011
`define JMP	1100	//RET
`define LEA	1110
`define TRAP 1111
